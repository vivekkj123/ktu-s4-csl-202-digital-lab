module OR_GATE(
	input A,
	input B,
	output Y
);

assign Y =  A||B;

endmodule;