module NOT_GATE(
	input A,
	output Y
);
assign Y = ~A;
endmodule;
